module processor(input clk);






endmodule
